module couter_circuit {
    input logic CLK, RST,
};