module top (
	input logic BTN0,
	output logic LED0_G
	);

	assign LED0_G = BTN0;

endmodule
